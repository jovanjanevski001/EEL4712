-- Jovan Janevski
-- UF-ID: 8591-9111
-- University of Florida

-- This tb tests the functionality of our 4-bit ripple carry adder

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity adder_tb is
end adder_tb;


architecture TB of adder_tb is 

signal input1, input2, sum : std_logic_vector(3 downto 0);
signal carry_in, carry_out : std_logic;

begin

	UUT: entity work.adder
		port map (
			input1		=>	input1,
			input2		=>	input2,
			carry_in	=>	carry_in,
			
			sum			=>	sum,
			carry_out	=>	carry_out
		);

	process
	
		-- function to check the sum
		function sum_check (
			in1, in2, c_in	:	integer)
			return std_logic_vector is
		begin 
			return std_logic_vector(to_unsigned((in1 + in2 + c_in) mod 16, 4));
		end sum_check;
		
		-- function to check carry_out
		function carry_out_check (
			in1, in2, c_in	:	integer)
			return std_logic is
		begin
			if (in1 + in2 + c_in > 15) then 
				return '1';
			else
				return '0';
			end if;
		end carry_out_check;
		
	begin 
		for i in 0 to 15 loop
			for j in 0 to 15 loop
				for k in 0 to 1 loop
					
					input1		<=	std_logic_vector(to_unsigned(i, 4));
					input2		<=	std_logic_vector(to_unsigned(j, 4));
					carry_in 	<= std_logic(to_unsigned(k, 1)(0));
					
					wait for 20 ns;
					assert(sum <= sum_check(i,j,k)) report "Incorrect Sum!" severity warning;
					assert(carry_out <= carry_out_check(i,j,k)) report "Incorrect Carry!" severity warning;

				end loop; -- k
			end loop; -- j
		end loop; -- i
		
		report "SIMULATION FINISHED!!!";
		wait;
	end process;
end TB;